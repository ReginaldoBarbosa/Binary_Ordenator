ENTITY teste_lab01 IS 
END ENTITY;

ARCHITECTURE simulacao OF teste_lab01 IS
	COMPONENT blocoFinal IS 
		PORT(A,B,C,D,E,F,G,H: IN bit; S1,S2,S3,S4,S5,S6,S7,S8: OUT bit);
	END COMPONENT;
	SIGNAL A,B,C,D,E,F,G,H,S1,S2,S3,S4,S5,S6,S7,S8: bit;
	
BEGIN

	tb: blocoFinal PORT MAP(A,B,C,D,E,F,G,H,S1,S2,S3,S4,S5,S6,S7,S8);
	PROCESS
		BEGIN
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 100 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 100 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 100 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 100 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 100 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 100 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 100 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '0'; E <= '0'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 100 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 100 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 100 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 100 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 100 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 100 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '0'; E <= '1'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '0'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '1'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '0'; D <= '1'; E <= '1'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 50 ns;	
		
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '0'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '0'; E <= '1'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 50 ns;	
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '0'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '0'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '0'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '0'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '0'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '1'; G <= '0'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '1'; G <= '0'; H <= '1'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '1'; G <= '1'; H <= '0'; WAIT FOR 50 ns;
			A <= '0'; B <= '0'; C <= '1'; D <= '1'; E <= '1'; F <= '1'; G <= '1'; H <= '1'; WAIT FOR 50 ns;
				
		END PROCESS;
END ARCHITECTURE; 
